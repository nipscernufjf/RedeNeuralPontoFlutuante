library verilog;
use verilog.vl_types.all;
entity teste_tb is
end teste_tb;
